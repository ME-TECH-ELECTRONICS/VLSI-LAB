module mux_4x1(y,s0,s1,d0,d1,d2,d3);
    input d0,d1,d2,d3,s0,s1;
    output y;
    wire ss_0
endmodule