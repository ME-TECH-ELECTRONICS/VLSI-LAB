class Payload;
    int payloadLen  = 1;
    rand bit[7:0] data;
    
endclass

class Header;

endclass