interface intf;
	logic a;
	logic b;
  	logic c;
endinterface