module dff ();
    
endmodule

module tb();
    clk=0;
    always #5 clk=~clk;
    initial begin
         
        
            
    end
    
endmodule