module array_types();
    int arr[3] = {20,40,34};
    string arr[3] {"Hello","World","!"};
    string arr3[];
    int arr4[string];
    
    
    endtask
    initial begin
        
        
    end
endmodule