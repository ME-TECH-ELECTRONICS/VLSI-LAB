module mux_4x1(y,s0,s1,d0,d1,d2,d3);
    input d0,d1,d2,d3,s0,s1;
    output y;
    wire s_0,s_1,t0,t1,t2,t3;
    and();
    and();
    and();
    and();
endmodule