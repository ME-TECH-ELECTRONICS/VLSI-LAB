class Scoreboard;
    mailbox scb_mbx;
    function new();
        
    endfunction 
endclass