interface dut_connector;
    logic[3:0] a;
    logic[3:0] b;
    logic[3:0] c;
endinterface