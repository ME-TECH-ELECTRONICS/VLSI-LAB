module tb ();
    int arr[] = {12,23,44};
    initial begin
        $display("%0d",arr[0]);
    end
endmodule