module partition_A (input wire N11, N130, N53, N380, N354, N373, N282, N345, N188, N376, N158, N105, N260, N122, N429, N276, N174, N267, N242, N285, N223, N17, N250, N415, N378, N356, N151, N432, N126, N186, N177, N142, N352, N418, N76, N343, N420, N134, N183, N336, N213, N1, N428, N60, N273, N404, N27, N421, N430, N292, N150, N348, N30, N243, N349, N146, N159, N425, N115, N251, N350, N393, N374, N375, N414, N47, N264, N147, N431, N360, N95, N259, N199, N108, N300, N305, N40, N381, N86, N184, N24, N351, N357, N355, N263, N377, N92, N82, N123, N191, N233, N224, N288, N8, N302, N330, N66, N4, N304, N196, N189, N258, N399, N338, N291, N190, N168, N379, N333, N89, N339, N257, N43, N340, N386, N256, N69, N422, N143, N307, N308, N230, N254, N289, N255, N370, N246, N411, N192, N139, N194, N342, N118, N347, N14, N334, N119, N157, N417, N73, N227, N37, N34, N239, N419, N306, N198, N332, N319, N247, N371, N63, N102, N165, N335, N372, N138, N127, N203, N301, N185, N99, N294, N193, N112, N50, N162, N341, N346, N195, N293, N296, N171, N131, N416, N21, N79, N197, N56, N180, N407, N309, N290, N187, N270, N353, N331, N279, N135, N154, N303, N236, N329, N295, N337, N344, output wire out);
    not     NOT1_1      (N118, N1, out);
    not     NOT1_2      (N119, N4, out);
    not     NOT1_3      (N122, N11, out);
    not     NOT1_4      (N123, N17, out);
    not     NOT1_9      (N134, N50, out);
    not     NOT1_10     (N135, N56, out);
    not     NOT1_13     (N142, N76, out);
    not     NOT1_16     (N147, N95, out);
    not     NOT1_17     (N150, N102, out);
    not     NOT1_18     (N151, N108, out);
    nand    NAND2_19    (N154, N118, N4, out);
    nor     NOR2_20     (N157, N8, N119, out);
    nor     NOR2_21     (N158, N14, N119, out);
    nand    NAND2_22    (N159, N122, N17, out);
    nand    NAND2_23    (N162, N126, N30, out);
    nand    NAND2_26    (N171, N138, N69, out);
    nand    NAND2_27    (N174, N142, N82, out);
    nand    NAND2_28    (N177, N146, N95, out);
    nand    NAND2_29    (N180, N150, N108, out);
    nor     NOR2_33     (N186, N40, N127, out);
    nor     NOR2_36     (N189, N60, N135, out);
    nor     NOR2_39     (N192, N79, N139, out);
    nor     NOR2_41     (N194, N92, N143, out);
    nor     NOR2_42     (N195, N99, N147, out);
    and     AND9_46     (N199, N154, N159, N162, N165, N168, N171, N174, N177, N180, out);
    not     NOT1_48     (N213, N199, out);
    xor     XOR2_53     (N233, N203, N165, out);
    xor     XOR2_54     (N236, N203, N168, out);
    xor     XOR2_57     (N243, N203, N174, out);
    nand    NAND2_58    (N246, N213, N11, out);
    nand    NAND2_60    (N250, N213, N24, out);
    nand    NAND2_62    (N254, N213, N37, out);
    nand    NAND2_63    (N255, N213, N50, out);
    nand    NAND2_64    (N256, N213, N63, out);
    nand    NAND2_67    (N259, N213, N102, out);
    nand    NAND2_68    (N260, N224, N157, out);
    nand    NAND2_70    (N264, N227, N183, out);
    nand    NAND2_72    (N270, N233, N187, out);
    nand    NAND2_74    (N276, N239, N191, out);
    nand    NAND2_75    (N279, N243, N193, out);
    nand    NAND2_77    (N285, N251, N197, out);
    nand    NAND2_78    (N288, N227, N184, out);
    nand    NAND2_80    (N290, N233, N188, out);
    nand    NAND2_83    (N293, N243, N194, out);
    nand    NAND2_84    (N294, N247, N196, out);
    nand    NAND2_85    (N295, N251, N198, out);
    and     AND9_86     (N296, N260, N264, N267, N270, N273, N276, N279, N282, N285, out);
    not     NOT1_87     (N300, N263, out);
    not     NOT1_93     (N306, N293, out);
    not     NOT1_94     (N307, N294, out);
    not     NOT1_96     (N309, N296, out);
    nand    NAND2_103   (N334, N8, N319, out);
    xor     XOR2_104    (N335, N309, N273, out);
    nand    NAND2_105   (N336, N319, N21, out);
    xor     XOR2_106    (N337, N309, N276, out);
    nand    NAND2_107   (N338, N319, N34, out);
    xor     XOR2_108    (N339, N309, N279, out);
    nand    NAND2_111   (N342, N319, N60, out);
    xor     XOR2_112    (N343, N309, N285, out);
    nand    NAND2_113   (N344, N319, N73, out);
    nand    NAND2_116   (N347, N319, N112, out);
    nand    NAND2_117   (N348, N330, N300, out);
    nand    NAND2_118   (N349, N331, N301, out);
    nand    NAND2_120   (N351, N333, N303, out);
    nand    NAND2_122   (N353, N337, N305, out);
    nand    NAND2_123   (N354, N339, N306, out);
    nand    NAND2_125   (N356, N343, N308, out);
    nand    NAND2_129   (N371, N14, N360, out);
    nand    NAND2_131   (N373, N360, N40, out);
    nand    NAND2_133   (N375, N360, N66, out);
    nand    NAND2_136   (N378, N360, N105, out);
    nand    NAND4_140   (N386, N250, N338, N373, N30, out);
    not     NOT1_147    (N415, N380, out);
    and     AND8_148    (N416, N381, N386, N393, N399, N404, N407, N411, N414, out);
    not     NOT1_149    (N417, N393, out);
    not     NOT1_151    (N419, N407, out);
    nand    NAND2_154   (N422, N386, N417, out);
    nand    NAND3_156   (N428, N399, N393, N419, out);
    nand    NAND4_158   (N430, N381, N386, N422, N399, out);
endmodule

module partition_B (input wire N11, N130, N53, N380, N354, N373, N282, N345, N188, N376, N158, N105, N260, N122, N429, N276, N174, N267, N242, N285, N223, N17, N250, N415, N378, N356, N151, N432, N126, N186, N177, N142, N352, N418, N76, N343, N420, N134, N183, N336, N213, N1, N428, N60, N273, N404, N27, N421, N430, N292, N150, N348, N30, N243, N349, N146, N159, N425, N115, N251, N350, N393, N374, N375, N414, N47, N264, N147, N431, N360, N95, N259, N199, N108, N300, N305, N40, N381, N86, N184, N24, N351, N357, N355, N263, N377, N92, N82, N123, N191, N233, N224, N288, N8, N302, N330, N66, N4, N304, N196, N189, N258, N399, N338, N291, N190, N168, N379, N333, N89, N339, N257, N43, N340, N386, N256, N69, N422, N143, N307, N308, N230, N254, N289, N255, N370, N246, N411, N192, N139, N194, N342, N118, N347, N14, N334, N119, N157, N417, N73, N227, N37, N34, N239, N419, N306, N198, N332, N319, N247, N371, N63, N102, N165, N335, N372, N138, N127, N203, N301, N185, N99, N294, N193, N112, N50, N162, N341, N346, N195, N293, N296, N171, N131, N416, N21, N79, N197, N56, N180, N407, N309, N290, N187, N270, N353, N331, N279, N135, N154, N303, N236, N329, N295, N337, N344, output wire out);
    not     NOT1_5      (N126, N24, out);
    not     NOT1_6      (N127, N30, out);
    not     NOT1_7      (N130, N37, out);
    not     NOT1_8      (N131, N43, out);
    not     NOT1_11     (N138, N63, out);
    not     NOT1_12     (N139, N69, out);
    not     NOT1_14     (N143, N82, out);
    not     NOT1_15     (N146, N89, out);
    nand    NAND2_24    (N165, N130, N43, out);
    nand    NAND2_25    (N168, N134, N56, out);
    nor     NOR2_30     (N183, N21, N123, out);
    nor     NOR2_31     (N184, N27, N123, out);
    nor     NOR2_32     (N185, N34, N127, out);
    nor     NOR2_34     (N187, N47, N131, out);
    nor     NOR2_35     (N188, N53, N131, out);
    nor     NOR2_37     (N190, N66, N135, out);
    nor     NOR2_38     (N191, N73, N139, out);
    nor     NOR2_40     (N193, N86, N143, out);
    nor     NOR2_43     (N196, N105, N147, out);
    nor     NOR2_44     (N197, N112, N151, out);
    nor     NOR2_45     (N198, N115, N151, out);
    not     NOT1_47     (N203, N199, out);
    not     NOT1_49     (N223, N199, out);
    xor     XOR2_50     (N224, N203, N154, out);
    xor     XOR2_51     (N227, N203, N159, out);
    xor     XOR2_52     (N230, N203, N162, out);
    xor     XOR2_55     (N239, N203, N171, out);
    nand    NAND2_56    (N242, N1, N213, out);
    xor     XOR2_59     (N247, N203, N177, out);
    xor     XOR2_61     (N251, N203, N180, out);
    nand    NAND2_65    (N257, N213, N76, out);
    nand    NAND2_66    (N258, N213, N89, out);
    nand    NAND2_69    (N263, N224, N158, out);
    nand    NAND2_71    (N267, N230, N185, out);
    nand    NAND2_73    (N273, N236, N189, out);
    nand    NAND2_76    (N282, N247, N195, out);
    nand    NAND2_79    (N289, N230, N186, out);
    nand    NAND2_81    (N291, N236, N190, out);
    nand    NAND2_82    (N292, N239, N192, out);
    not     NOT1_88     (N301, N288, out);
    not     NOT1_89     (N302, N289, out);
    not     NOT1_90     (N303, N290, out);
    not     NOT1_91     (N304, N291, out);
    not     NOT1_92     (N305, N292, out);
    not     NOT1_95     (N308, N295, out);
    not     NOT1_97     (N319, N296, out);
    not     NOT1_98     (N329, N296, out);
    xor     XOR2_99     (N330, N309, N260, out);
    xor     XOR2_100    (N331, N309, N264, out);
    xor     XOR2_101    (N332, N309, N267, out);
    xor     XOR2_102    (N333, N309, N270, out);
    nand    NAND2_109   (N340, N319, N47, out);
    xor     XOR2_110    (N341, N309, N282, out);
    nand    NAND2_114   (N345, N319, N86, out);
    nand    NAND2_115   (N346, N319, N99, out);
    nand    NAND2_119   (N350, N332, N302, out);
    nand    NAND2_121   (N352, N335, N304, out);
    nand    NAND2_124   (N355, N341, N307, out);
    and     AND9_126    (N357, N348, N349, N350, N351, N352, N353, N354, N355, N356, out);
    not     NOT1_127    (N360, N357, out);
    not     NOT1_128    (N370, N357, out);
    nand    NAND2_130   (N372, N360, N27, out);
    nand    NAND2_132   (N374, N360, N53, out);
    nand    NAND2_134   (N376, N360, N79, out);
    nand    NAND2_135   (N377, N360, N92, out);
    nand    NAND2_137   (N379, N360, N115, out);
    nand    NAND4_138   (N380, N4, N242, N334, N371, out);
    nand    NAND4_139   (N381, N246, N336, N372, N17, out);
    nand    NAND4_141   (N393, N254, N340, N374, N43, out);
    nand    NAND4_142   (N399, N255, N342, N375, N56, out);
    nand    NAND4_143   (N404, N256, N344, N376, N69, out);
    nand    NAND4_144   (N407, N257, N345, N377, N82, out);
    nand    NAND4_145   (N411, N258, N346, N378, N95, out);
    nand    NAND4_146   (N414, N259, N347, N379, N108, out);
    not     NOT1_150    (N418, N404, out);
    not     NOT1_152    (N420, N411, out);
    nor     NOR2_153    (N421, N415, N416, out);
    nand    NAND4_155   (N425, N386, N393, N418, N399, out);
    nand    NAND4_157   (N429, N386, N393, N407, N420, out);
    nand    NAND4_159   (N431, N381, N386, N425, N428, out);
    nand    NAND4_160   (N432, N381, N422, N425, N429, out);
endmodule


module full_circuit(input wire N11, N130, N53, N380, N354, N373, N282, N345, N188, N376, N158, N105, N260, N122, N429, N276, N174, N267, N242, N285, N223, N17, N250, N415, N378, N356, N151, N432, N126, N186, N177, N142, N352, N418, N76, N343, N420, N134, N183, N336, N213, N1, N428, N60, N273, N404, N27, N421, N430, N292, N150, N348, N30, N243, N349, N146, N159, N425, N115, N251, N350, N393, N374, N375, N414, N47, N264, N147, N431, N360, N95, N259, N199, N108, N300, N305, N40, N381, N86, N184, N24, N351, N357, N355, N263, N377, N92, N82, N123, N191, N233, N224, N288, N8, N302, N330, N66, N4, N304, N196, N189, N258, N399, N338, N291, N190, N168, N379, N333, N89, N339, N257, N43, N340, N386, N256, N69, N422, N143, N307, N308, N230, N254, N289, N255, N370, N246, N411, N192, N139, N194, N342, N118, N347, N14, N334, N119, N157, N417, N73, N227, N37, N34, N239, N419, N306, N198, N332, N319, N247, N371, N63, N102, N165, N335, N372, N138, N127, N203, N301, N185, N99, N294, N193, N112, N50, N162, N341, N346, N195, N293, N296, N171, N131, N416, N21, N79, N197, N56, N180, N407, N309, N290, N187, N270, N353, N331, N279, N135, N154, N303, N236, N329, N295, N337, N344, output wire out);
    wire mid;
    partition_A A (N11, N130, N53, N380, N354, N373, N282, N345, N188, N376, N158, N105, N260, N122, N429, N276, N174, N267, N242, N285, N223, N17, N250, N415, N378, N356, N151, N432, N126, N186, N177, N142, N352, N418, N76, N343, N420, N134, N183, N336, N213, N1, N428, N60, N273, N404, N27, N421, N430, N292, N150, N348, N30, N243, N349, N146, N159, N425, N115, N251, N350, N393, N374, N375, N414, N47, N264, N147, N431, N360, N95, N259, N199, N108, N300, N305, N40, N381, N86, N184, N24, N351, N357, N355, N263, N377, N92, N82, N123, N191, N233, N224, N288, N8, N302, N330, N66, N4, N304, N196, N189, N258, N399, N338, N291, N190, N168, N379, N333, N89, N339, N257, N43, N340, N386, N256, N69, N422, N143, N307, N308, N230, N254, N289, N255, N370, N246, N411, N192, N139, N194, N342, N118, N347, N14, N334, N119, N157, N417, N73, N227, N37, N34, N239, N419, N306, N198, N332, N319, N247, N371, N63, N102, N165, N335, N372, N138, N127, N203, N301, N185, N99, N294, N193, N112, N50, N162, N341, N346, N195, N293, N296, N171, N131, N416, N21, N79, N197, N56, N180, N407, N309, N290, N187, N270, N353, N331, N279, N135, N154, N303, N236, N329, N295, N337, N344, mid);
    partition_B B (N11, N130, N53, N380, N354, N373, N282, N345, N188, N376, N158, N105, N260, N122, N429, N276, N174, N267, N242, N285, N223, N17, N250, N415, N378, N356, N151, N432, N126, N186, N177, N142, N352, N418, N76, N343, N420, N134, N183, N336, N213, N1, N428, N60, N273, N404, N27, N421, N430, N292, N150, N348, N30, N243, N349, N146, N159, N425, N115, N251, N350, N393, N374, N375, N414, N47, N264, N147, N431, N360, N95, N259, N199, N108, N300, N305, N40, N381, N86, N184, N24, N351, N357, N355, N263, N377, N92, N82, N123, N191, N233, N224, N288, N8, N302, N330, N66, N4, N304, N196, N189, N258, N399, N338, N291, N190, N168, N379, N333, N89, N339, N257, N43, N340, N386, N256, N69, N422, N143, N307, N308, N230, N254, N289, N255, N370, N246, N411, N192, N139, N194, N342, N118, N347, N14, N334, N119, N157, N417, N73, N227, N37, N34, N239, N419, N306, N198, N332, N319, N247, N371, N63, N102, N165, N335, N372, N138, N127, N203, N301, N185, N99, N294, N193, N112, N50, N162, N341, N346, N195, N293, N296, N171, N131, N416, N21, N79, N197, N56, N180, N407, N309, N290, N187, N270, N353, N331, N279, N135, N154, N303, N236, N329, N295, N337, N344, out);
endmodule
    

    

module testbench;

    reg N11, N130, N53, N380, N354, N373, N282, N345, N188, N376, N158, N105, N260, N122, N429, N276, N174, N267, N242, N285, N223, N17, N250, N415, N378, N356, N151, N432, N126, N186, N177, N142, N352, N418, N76, N343, N420, N134, N183, N336, N213, N1, N428, N60, N273, N404, N27, N421, N430, N292, N150, N348, N30, N243, N349, N146, N159, N425, N115, N251, N350, N393, N374, N375, N414, N47, N264, N147, N431, N360, N95, N259, N199, N108, N300, N305, N40, N381, N86, N184, N24, N351, N357, N355, N263, N377, N92, N82, N123, N191, N233, N224, N288, N8, N302, N330, N66, N4, N304, N196, N189, N258, N399, N338, N291, N190, N168, N379, N333, N89, N339, N257, N43, N340, N386, N256, N69, N422, N143, N307, N308, N230, N254, N289, N255, N370, N246, N411, N192, N139, N194, N342, N118, N347, N14, N334, N119, N157, N417, N73, N227, N37, N34, N239, N419, N306, N198, N332, N319, N247, N371, N63, N102, N165, N335, N372, N138, N127, N203, N301, N185, N99, N294, N193, N112, N50, N162, N341, N346, N195, N293, N296, N171, N131, N416, N21, N79, N197, N56, N180, N407, N309, N290, N187, N270, N353, N331, N279, N135, N154, N303, N236, N329, N295, N337, N344;
    wire out;
    full_circuit uut (N11, N130, N53, N380, N354, N373, N282, N345, N188, N376, N158, N105, N260, N122, N429, N276, N174, N267, N242, N285, N223, N17, N250, N415, N378, N356, N151, N432, N126, N186, N177, N142, N352, N418, N76, N343, N420, N134, N183, N336, N213, N1, N428, N60, N273, N404, N27, N421, N430, N292, N150, N348, N30, N243, N349, N146, N159, N425, N115, N251, N350, N393, N374, N375, N414, N47, N264, N147, N431, N360, N95, N259, N199, N108, N300, N305, N40, N381, N86, N184, N24, N351, N357, N355, N263, N377, N92, N82, N123, N191, N233, N224, N288, N8, N302, N330, N66, N4, N304, N196, N189, N258, N399, N338, N291, N190, N168, N379, N333, N89, N339, N257, N43, N340, N386, N256, N69, N422, N143, N307, N308, N230, N254, N289, N255, N370, N246, N411, N192, N139, N194, N342, N118, N347, N14, N334, N119, N157, N417, N73, N227, N37, N34, N239, N419, N306, N198, N332, N319, N247, N371, N63, N102, N165, N335, N372, N138, N127, N203, N301, N185, N99, N294, N193, N112, N50, N162, N341, N346, N195, N293, N296, N171, N131, N416, N21, N79, N197, N56, N180, N407, N309, N290, N187, N270, N353, N331, N279, N135, N154, N303, N236, N329, N295, N337, N344, out);

    initial begin
        $dumpfile("c432_tb.vcd");
        $dumpvars(0, testbench);
        $monitor("Time=%0t | Output: %b", $time, out);
        N11     = 1'b0;
        N130    = 1'b0;
        N53     = 1'b0;
        N380    = 1'b0;
        N354    = 1'b0;
        N373    = 1'b0;
        N282    = 1'b0;
        N345    = 1'b0;
        N188    = 1'b0;
        N376    = 1'b0;
        N158    = 1'b0;
        N105    = 1'b0;
        N260    = 1'b0;
        N122    = 1'b0;
        N429    = 1'b0;
        N276    = 1'b0;
        N174    = 1'b0;
        N267    = 1'b0;
        N242    = 1'b0;
        N285    = 1'b0;
        N223    = 1'b0;
        N17     = 1'b0;
        N250    = 1'b0;
        N415    = 1'b0;
        N378    = 1'b0;
        N356    = 1'b0;
        N151    = 1'b0;
        N432    = 1'b0;
        N126    = 1'b0;
        N186    = 1'b0;
        N177    = 1'b0;
        N142    = 1'b0;
        N352    = 1'b0;
        N418    = 1'b0;
        N76     = 1'b0;
        N343    = 1'b0;
        N420    = 1'b0;
        N134    = 1'b0;
        N183    = 1'b0;
        N336    = 1'b0;
        N213    = 1'b0;
        N1      = 1'b0;
        N428    = 1'b0;
        N60     = 1'b0;
        N273    = 1'b0;
        N404    = 1'b0;
        N27     = 1'b0;
        N421    = 1'b0;
        N430    = 1'b0;
        N292    = 1'b0;
        N150    = 1'b0;
        N348    = 1'b0;
        N30     = 1'b0;
        N243    = 1'b0;
        N349    = 1'b0;
        N146    = 1'b0;
        N159    = 1'b0;
        N425    = 1'b0;
        N115    = 1'b0;
        N251    = 1'b0;
        N350    = 1'b0;
        N393    = 1'b0;
        N374    = 1'b0;
        N375    = 1'b0;
        N414    = 1'b0;
        N47     = 1'b0;
        N264    = 1'b0;
        N147    = 1'b0;
        N431    = 1'b0;
        N360    = 1'b0;
        N95     = 1'b0;
        N259    = 1'b0;
        N199    = 1'b0;
        N108    = 1'b0;
        N300    = 1'b0;
        N305    = 1'b0;
        N40     = 1'b0;
        N381    = 1'b0;
        N86     = 1'b0;
        N184    = 1'b0;
        N24     = 1'b0;
        N351    = 1'b0;
        N357    = 1'b0;
        N355    = 1'b0;
        N263    = 1'b0;
        N377    = 1'b0;
        N92     = 1'b0;
        N82     = 1'b0;
        N123    = 1'b0;
        N191    = 1'b0;
        N233    = 1'b0;
        N224    = 1'b0;
        N288    = 1'b0;
        N8      = 1'b0;
        N302    = 1'b0;
        N330    = 1'b0;
        N66     = 1'b0;
        N4      = 1'b0;
        N304    = 1'b0;
        N196    = 1'b0;
        N189    = 1'b0;
        N258    = 1'b0;
        N399    = 1'b0;
        N338    = 1'b0;
        N291    = 1'b0;
        N190    = 1'b0;
        N168    = 1'b0;
        N379    = 1'b0;
        N333    = 1'b0;
        N89     = 1'b0;
        N339    = 1'b0;
        N257    = 1'b0;
        N43     = 1'b0;
        N340    = 1'b0;
        N386    = 1'b0;
        N256    = 1'b0;
        N69     = 1'b0;
        N422    = 1'b0;
        N143    = 1'b0;
        N307    = 1'b0;
        N308    = 1'b0;
        N230    = 1'b0;
        N254    = 1'b0;
        N289    = 1'b0;
        N255    = 1'b0;
        N370    = 1'b0;
        N246    = 1'b0;
        N411    = 1'b0;
        N192    = 1'b0;
        N139    = 1'b0;
        N194    = 1'b0;
        N342    = 1'b0;
        N118    = 1'b0;
        N347    = 1'b0;
        N14     = 1'b0;
        N334    = 1'b0;
        N119    = 1'b0;
        N157    = 1'b0;
        N417    = 1'b0;
        N73     = 1'b0;
        N227    = 1'b0;
        N37     = 1'b0;
        N34     = 1'b0;
        N239    = 1'b0;
        N419    = 1'b0;
        N306    = 1'b0;
        N198    = 1'b0;
        N332    = 1'b0;
        N319    = 1'b0;
        N247    = 1'b0;
        N371    = 1'b0;
        N63     = 1'b0;
        N102    = 1'b0;
        N165    = 1'b0;
        N335    = 1'b0;
        N372    = 1'b0;
        N138    = 1'b0;
        N127    = 1'b0;
        N203    = 1'b0;
        N301    = 1'b0;
        N185    = 1'b0;
        N99     = 1'b0;
        N294    = 1'b0;
        N193    = 1'b0;
        N112    = 1'b0;
        N50     = 1'b0;
        N162    = 1'b0;
        N341    = 1'b0;
        N346    = 1'b0;
        N195    = 1'b0;
        N293    = 1'b0;
        N296    = 1'b0;
        N171    = 1'b0;
        N131    = 1'b0;
        N416    = 1'b0;
        N21     = 1'b0;
        N79     = 1'b0;
        N197    = 1'b0;
        N56     = 1'b0;
        N180    = 1'b0;
        N407    = 1'b0;
        N309    = 1'b0;
        N290    = 1'b0;
        N187    = 1'b0;
        N270    = 1'b0;
        N353    = 1'b0;
        N331    = 1'b0;
        N279    = 1'b0;
        N135    = 1'b0;
        N154    = 1'b0;
        N303    = 1'b0;
        N236    = 1'b0;
        N329    = 1'b0;
        N295    = 1'b0;
        N337    = 1'b0;
        N344    = 1'b0;;
        #10;
        N11     = $random; #10;
        N130    = $random; #10;
        N53     = $random; #10;
        N380    = $random; #10;
        N354    = $random; #10;
        N373    = $random; #10;
        N282    = $random; #10;
        N345    = $random; #10;
        N188    = $random; #10;
        N376    = $random; #10;
        N158    = $random; #10;
        N105    = $random; #10;
        N260    = $random; #10;
        N122    = $random; #10;
        N429    = $random; #10;
        N276    = $random; #10;
        N174    = $random; #10;
        N267    = $random; #10;
        N242    = $random; #10;
        N285    = $random; #10;
        N223    = $random; #10;
        N17     = $random; #10;
        N250    = $random; #10;
        N415    = $random; #10;
        N378    = $random; #10;
        N356    = $random; #10;
        N151    = $random; #10;
        N432    = $random; #10;
        N126    = $random; #10;
        N186    = $random; #10;
        N177    = $random; #10;
        N142    = $random; #10;
        N352    = $random; #10;
        N418    = $random; #10;
        N76     = $random; #10;
        N343    = $random; #10;
        N420    = $random; #10;
        N134    = $random; #10;
        N183    = $random; #10;
        N336    = $random; #10;
        N213    = $random; #10;
        N1      = $random; #10;
        N428    = $random; #10;
        N60     = $random; #10;
        N273    = $random; #10;
        N404    = $random; #10;
        N27     = $random; #10;
        N421    = $random; #10;
        N430    = $random; #10;
        N292    = $random; #10;
        N150    = $random; #10;
        N348    = $random; #10;
        N30     = $random; #10;
        N243    = $random; #10;
        N349    = $random; #10;
        N146    = $random; #10;
        N159    = $random; #10;
        N425    = $random; #10;
        N115    = $random; #10;
        N251    = $random; #10;
        N350    = $random; #10;
        N393    = $random; #10;
        N374    = $random; #10;
        N375    = $random; #10;
        N414    = $random; #10;
        N47     = $random; #10;
        N264    = $random; #10;
        N147    = $random; #10;
        N431    = $random; #10;
        N360    = $random; #10;
        N95     = $random; #10;
        N259    = $random; #10;
        N199    = $random; #10;
        N108    = $random; #10;
        N300    = $random; #10;
        N305    = $random; #10;
        N40     = $random; #10;
        N381    = $random; #10;
        N86     = $random; #10;
        N184    = $random; #10;
        N24     = $random; #10;
        N351    = $random; #10;
        N357    = $random; #10;
        N355    = $random; #10;
        N263    = $random; #10;
        N377    = $random; #10;
        N92     = $random; #10;
        N82     = $random; #10;
        N123    = $random; #10;
        N191    = $random; #10;
        N233    = $random; #10;
        N224    = $random; #10;
        N288    = $random; #10;
        N8      = $random; #10;
        N302    = $random; #10;
        N330    = $random; #10;
        N66     = $random; #10;
        N4      = $random; #10;
        N304    = $random; #10;
        N196    = $random; #10;
        N189    = $random; #10;
        N258    = $random; #10;
        N399    = $random; #10;
        N338    = $random; #10;
        N291    = $random; #10;
        N190    = $random; #10;
        N168    = $random; #10;
        N379    = $random; #10;
        N333    = $random; #10;
        N89     = $random; #10;
        N339    = $random; #10;
        N257    = $random; #10;
        N43     = $random; #10;
        N340    = $random; #10;
        N386    = $random; #10;
        N256    = $random; #10;
        N69     = $random; #10;
        N422    = $random; #10;
        N143    = $random; #10;
        N307    = $random; #10;
        N308    = $random; #10;
        N230    = $random; #10;
        N254    = $random; #10;
        N289    = $random; #10;
        N255    = $random; #10;
        N370    = $random; #10;
        N246    = $random; #10;
        N411    = $random; #10;
        N192    = $random; #10;
        N139    = $random; #10;
        N194    = $random; #10;
        N342    = $random; #10;
        N118    = $random; #10;
        N347    = $random; #10;
        N14     = $random; #10;
        N334    = $random; #10;
        N119    = $random; #10;
        N157    = $random; #10;
        N417    = $random; #10;
        N73     = $random; #10;
        N227    = $random; #10;
        N37     = $random; #10;
        N34     = $random; #10;
        N239    = $random; #10;
        N419    = $random; #10;
        N306    = $random; #10;
        N198    = $random; #10;
        N332    = $random; #10;
        N319    = $random; #10;
        N247    = $random; #10;
        N371    = $random; #10;
        N63     = $random; #10;
        N102    = $random; #10;
        N165    = $random; #10;
        N335    = $random; #10;
        N372    = $random; #10;
        N138    = $random; #10;
        N127    = $random; #10;
        N203    = $random; #10;
        N301    = $random; #10;
        N185    = $random; #10;
        N99     = $random; #10;
        N294    = $random; #10;
        N193    = $random; #10;
        N112    = $random; #10;
        N50     = $random; #10;
        N162    = $random; #10;
        N341    = $random; #10;
        N346    = $random; #10;
        N195    = $random; #10;
        N293    = $random; #10;
        N296    = $random; #10;
        N171    = $random; #10;
        N131    = $random; #10;
        N416    = $random; #10;
        N21     = $random; #10;
        N79     = $random; #10;
        N197    = $random; #10;
        N56     = $random; #10;
        N180    = $random; #10;
        N407    = $random; #10;
        N309    = $random; #10;
        N290    = $random; #10;
        N187    = $random; #10;
        N270    = $random; #10;
        N353    = $random; #10;
        N331    = $random; #10;
        N279    = $random; #10;
        N135    = $random; #10;
        N154    = $random; #10;
        N303    = $random; #10;
        N236    = $random; #10;
        N329    = $random; #10;
        N295    = $random; #10;
        N337    = $random; #10;
        N344    = $random; #10;;
        #100;
        
        $finish;
    end

endmodule
    