module name ();
int array_types[4]={20,10,30};


end