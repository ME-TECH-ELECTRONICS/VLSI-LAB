class
module tb ();
    
endmodule