interface dut_connector;
    
endinterface