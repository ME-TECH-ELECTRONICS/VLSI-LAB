interface adder_intf();
    logic[7;0] a;
    logic[7;0] b;
    bit[7:0] sum;
    bit carry;
endinterface