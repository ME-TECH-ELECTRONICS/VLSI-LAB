interface adder_intf();
    logic a;
    logic b;
    logic c;
    bit sum;
    bit carry;
endinterface