`include "slave.sv"
`include "master.sv"

module apb_top(
  input logic PCLK, RST_N, TX, APB_SWRITE,
  input logic [8:0] APB_SLV_PADDR,
  input logic [7:0] APB_PWDATA,
  output logic [7:0] APB_PRDATA
);
  logic [7:0]PWDATA,PRDATA,PRDATA1,PRDATA2;
  logic [8:0]PADDR;         
  logic PREADY,PREADY1,PREADY2,PENABLE,PSEL1,PSEL2,PWRITE;
  
  assign PREADY = PADDR[8] ? PREADY2 : PREADY1 ;
  assign PRDATA = APB_SWRITE ? (PADDR[8] ? PRDATA2 : PRDATA1) : 8'dx ;
  
  APB_MASTER dut (CLK,RST_N,PREADY,PSLVERR,PRDATA,APB_SLV_PADDR,APB_PWDATA,TX,APB_SWRITE,PSEL1,PSEL2,PEN,PWRITE,PADDR,PWDATA, APB_PRDATA );

  APB_SLAVE slv1(CLK,RST_N,PWRITE,PSEL1,PEN,PADDR[7:0],PWDATA,PREADY1,PSLVERR,PRDATA1);
  APB_SLAVE slv2(CLK,RST_N,PWRITE,PSEL2,PEN,PADDR[7:0],PWDATA,PREADY2,PSLVERR,PRDATA2);
endmodule
