module APB_master (
    input wire clk,
    input wire rst,
    input wire pready,
    input wire [31:0] prdata,
    output reg psel,
    output reg pen,
    output reg pwr,
    output reg pslverr,
    output reg [31:0] pwdata,
    output reg [31:0] pwdata,
);
    
endmodule