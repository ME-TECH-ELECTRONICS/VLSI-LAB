class first;
    int data = 10;
    function first copy();
        copy = new();
        copy.data = data;
    endfunction 
endclass 

class second;
    function new();
        
    endfunction 
endclass 