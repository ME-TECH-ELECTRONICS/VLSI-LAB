module SPI_PERIFERIAL (
    ports
);
    
endmodule