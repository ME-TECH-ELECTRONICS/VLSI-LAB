module tb ();
    int arr[5];
    
endmodule